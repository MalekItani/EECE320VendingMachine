library ieee;
use ieee.std_logic_1164.all;
entity itemToPrice is
  port (
    itemNumber: in std_logic_vector(11 downto 0);
    price: out std_logic_vector(4 downto 0)
  );
end entity;

architecture archItemToPrice of ItemToPrice is
begin
  with itemNumber
  select price <= "00010" when "001000000010" | "001000000011" | "001000000101" | "001000000110" | -- 202, 203, 205, 206
                               "001100000001" | "010000001000" | "010000001011" | "010000010010", -- 301, 408, 411, 412
                  "00100" when "000100000001" | "000100000010" | "000100000011" | "001000000001" |-- 101, 102, 103, 201
                               "001100000010" | "001100000110" | "010000000111" | "010000001001" | "010000010000" | -- 302, 306, 407, 409, 410
                               "011000000001" | "011000000010" | "011000000011" | "011000000100" | "011000000101" | -- 601 - 605
                               "011000000110" | "011000000111" | "011000001000" | "011000001001" | "011000010000", -- 606 - 610 XX
                  "00110" when "000100000100" | "000100000101" | "000100000110" | "001000000100" |-- 104, 105, 106, 204
                               "001100000100" | "001100000101" | "010000000001" | "010000000010" | "010000000011" | "010000000100" |-- 304, 305, 401, 402, 403, 404
                               "010100000001" | "010100000010" | "010100000011" | "010100000100", -- 501, 502, 503, 504
                  "01000" when "001100000011" | "010000000101" | "010000000110" | "010100000101" | "010100000110" | "010100000111",-- 303, 405, 406, 505, 506, 507
                  "01100" when "010100001000" | "010100001001", -- 508, 509,
                  "01110" when "010100010000", -- 510
                  "00000" when others;

end architecture;
