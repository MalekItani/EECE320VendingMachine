library ieee;
use ieee.std_logic_1164.all;
entity itemToPrice is
  port (
    itemNumber: in std_logic_vector(9 downto 0);
    price: out std_logic_vector(4 downto 0)
  );
end entity;

architecture archItemToPrice of ItemToPrice is
begin
  with itemNumber
  select price <= "00010" when "0011001010" | "0011001011" | "0011001101" | "0011001110" | -- 202, 203, 205, 206
                               "0100101101" | "0110011000" | "0110011011" | "0110011100", -- 301, 408, 411, 412
                  "00100" when "0001100101" | "0001100110" | "0001100111" | "0011001001" |-- 101, 102, 103, 201
                               "0100101110" | "0100110010" | "0110010111" | "0110011001" | "0110011010" | -- 302, 306, 407, 409, 410
                               "1001011001" | "1001011010" | "1001011011" | "1001011100" | "1001011101" | -- 601 - 605
                               "1001011110" | "1001011111" | "1001100000" | "1001100001" | "1001100010", -- 606 - 610
                  "00110" when "0001101000" | "0001101001" | "0001101010" | "0011001100" |-- 104, 105, 106, 204
                               "0100110000" | "0100110001" | "0110010001" | "0110010010" | "0110010011" | "0110010100" |-- 304, 305, 401, 402, 403, 404
                               "0111110101" | "0111110110" | "0111110111" | "0111111000", -- 501, 502, 503, 504
                  "01000" when "0100101111" | "0110010101" | "0110010110" | "0111111001" | "0111111010" | "0111111011",-- 303, 405, 406, 505, 506, 507
                  "01100" when "0111111100" | "0111111101", -- 508, 509,
                  "01110" when "0111111110", -- 510
                  "11111" when others;

end architecture;
